module ysyx_22041211_branchJmp #(parameter DATA_LEN = 32)(
	input		                		zero,
	input		                        branch,
	input 		                        jmp,
	output		                        PCSrc
);
    assign PCSrc = jmp | (zero & branch);

endmodule