module ysyx_22041211_branchJmp(
	input		                		zero,
	input		                        branch,
	input 		                        jmp,
	output		  [1:0]                 PCSrc
);
    //00--default
    //01
    //10

endmodule

